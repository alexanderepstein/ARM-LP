module PC(output reg[31:0] readAddress);

endmodule 
