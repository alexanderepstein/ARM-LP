module Controller(input[31:0] address, output wire reg2Loc,
    output wire unconditionalBranch, output wire branch, output wire memRead,
    output wire memToReg, output wire aluOP, output wire memWrite,
    output wire aluSRC, output wire regWrite, output reg [4:0] readRegister1,
    output reg [4:0] readRegister2, output reg [4:0] writeRegister) ;
    
    //Those only did the straight control

endmodule 