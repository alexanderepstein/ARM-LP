module OperationPrep(input wire regWrite, input [4:0] reg1, input[4:0] reg2,
 input[4:0] writeRegister, input[31:0] writeData, output reg [4:0] readData1,
 output reg[4:0] readData2, input wire aluSRC);

endmodule 
