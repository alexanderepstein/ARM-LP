module Controller() ;

endmodule 