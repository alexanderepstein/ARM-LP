module InstructionCache(input[31:0] address, output reg[31:0] instruction);

endmodule 