module DataCache();

endmodule 