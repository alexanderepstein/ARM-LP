module DataCache(input wire memWrite, input wire memRead, input wire memToReg,
 input[31:0] address, input[31:0] writeData, output reg [31:0] readData, input reg clock);

endmodule 
