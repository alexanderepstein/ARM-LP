module top();

endmodule 