module InstructionCache(input[31:0] address, output reg[31:0] instruction,
 input clock);

 	always @(posedge clock) begin

    end
endmodule 