module InstructionCache();

endmodule 