module Controller(input[31:0] address, output reg reg2LocOut,
    output reg unconditionalBranch, output reg branch, output reg memRead,
    output reg memToReg, output reg aluOP, output reg memWrite,
    output reg aluSRC, output reg regWrite, output reg [4:0] readRegister1,
    output reg [4:0] readRegister2, output reg [4:0] writeRegister,
    input wire reg2LocIn) ;
    
endmodule 