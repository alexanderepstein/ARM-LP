module DataCache(input wire memWrite, input wire memRead, input wire memToReg,
 input[31:0] address, input[3:0] writeData, output reg [31:0] readData, input clock);

endmodule 