module OperationPrep();

endmodule 