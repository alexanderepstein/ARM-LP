module PC();

endmodule 